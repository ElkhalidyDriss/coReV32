---------------------------------------------------------------------------------------
--  Author: Driss Elkhalidy , an embedded systems engineering student                -- 
--          at National Institute of Posts and Telecommunications , Rabat , Morocco. --
--  Description : Implementation of the top level entity for the coReV32.            --
--  Dependencies : rv_regFile.vhd ,rv_alu.vhd 
---------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity rv_core is 
end entity;


architecture rv_core_arch of rv_core is 


begin


end architecture;
